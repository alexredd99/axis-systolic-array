`define WK                  8        
`define WX                  8
`define WA                  32
`define WY                  32
`define LM                  1
`define LA                  1
`define AXI_WIDTH           128
`define AXI_ID_WIDTH        6
`define AXI_STRB_WIDTH      `AXI_WIDTH/8
`define AXI_MAX_BURST_LEN   32
`define AXI_ADDR_WIDTH	    32
`define AXIL_WIDTH          32
`define AXIL_ADDR_WIDTH     40
`define STRB_WIDTH          4 
`define AXIL_BASE_ADDR      32'hA0000000